`ifndef _%N_%E_INCLUDED
`define _%N_%E_INCLUDED

/** @file */

`include "%n.svh"

%@

`endif
