//------------------------------------------------------------------------------
//  Copyright (c) %Y Cisco Systems Inc. All rights reserved.
//  This software product contains the unpublished source code of
//  Cisco Systems Inc. The copyright notices above do not evidence
//  any actual or intended publication of such source code.
//
//  File Name:         %b
//
//  Language:          System Verilog
//
//  File Description:  %@
//
//  Initial Version:   %d %M %Y  By: %u
//
//------------------------------------------------------------------------------
//
// $Id: $

`include "%n.svh"
