// Copyright (C) Microsoft Corporation. All rights reserved.

`ifndef %N
`define %N

%@

`endif
