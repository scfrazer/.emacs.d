/** @file */

`include "%n.svh"

%@
