//--------------------------------------------------------------------------
//  Cisco Systems Inc.
//
//  Copyright (c) %Y Cisco Systems Inc.
//  All rights reserved
//
//  This software product contains the unpublished source code of
//  Cisco Systems Inc.
//
//  The copyright notices above do not evidence any actual or
//  intended publication of such source code.
//
//  File Name:          %b
//
//  Language:           SystemVerilog
//
//  File Description:   %[Description: %]
//
//  Initial Version:    %d %M %Y    By: %u
//
//--------------------------------------------------------------------------

/** @file */

`include "%n.svh"

%@