// Copyright (C) Microsoft Corporation. All rights reserved.
