// ----------------------------------------------------------------------------
//
//   Title    : %[Title: %]
//   Filename : %b
//   Language : SystemVerilog
//   Author   : %u
//
//   Description : %1
//
// ----------------------------------------------------------------------------
// Copyright (c) %Y by Cisco Systems, Inc
// This model is the confidential and proprietary property of Cisco and the
// possession or use of this file requires written permission from Cisco.
// ----------------------------------------------------------------------------

/** @file */

`include "%n.h"

%@
